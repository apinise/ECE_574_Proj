module fir_tb (
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic clk;
logic reset;

logic start;
logic done;

logic [11:0]  din;
logic [11:0]  dout;

logic [11:0]  chkDout;
logic 	      testbench_pass;
integer       fvectors, r;

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

fir_transpose DUT(
  .Clk(clk),
  .Hlt(reset),
  .Din(din),
  .Dout(dout)
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

initial begin
  fvectors = $fopen("../refC/vectors.txt", "r");
  if (fvectors == 0) begin
     $display("Could not open refC/vectors.txt");
     $finish;
  end
  
	clk = 0;
	din = 0;
	start = 0;
	testbench_pass = 1;
  
	reset = 1;
	@(posedge clk);
  #7;
  @(posedge clk);
	reset = 0;
  
	while (!$feof(fvectors))
	  begin
	     r = $fscanf(fvectors,"%d %d\n", din, chkDout);
       
	     @(posedge clk);
       
       $display("Din %d Dout %d chkDout %d OK %b", din, dout, chkDout, (dout == chkDout));
	     testbench_pass = testbench_pass && (dout == chkDout);	     
	  end

	$fclose(fvectors);
  
	if (testbench_pass)
	  $display("TESTBENCH PASSES");
	else
	  $display("TESTBENCH FAILS");
    
  $finish;
  
end

always begin
 #5 clk = ~clk;
end

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

endmodule