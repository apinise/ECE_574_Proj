/opt/cadence/libraries/gsclib045_all_v4.7/gsclib045/lef/gsclib045_macro.lef